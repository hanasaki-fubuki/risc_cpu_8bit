LIBRARY IEEE ;
USE IEEE.STD_LOGIC_1164.ALL ;
ENTITY REG8 IS 
	PORT (CLK : IN STD_LOGIC ;
	D : IN STD_LOGIC_VECTOR(7 DOWNTO 0) ;
	Q : OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END;
ARCHITECTURE bhv OF REG8 IS
	SIGNAL Q1 : STD_LOGIC_VECTOR(7 DOWNTO 0) ;
		BEGIN
			PROCESS (CLK,Q1)
				BEGIN
					IF CLK'EVENT AND CLK='1'
						THEN Q1<=d;
					END IF;
				END PROCESS;
			Q<=Q1;
		END bhv;
	